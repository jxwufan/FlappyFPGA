
 
 
 




window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"


      waveform add -signals /ret_back_tb/status
      waveform add -signals /ret_back_tb/ret_back_synth_inst/bmg_port/CLKA
      waveform add -signals /ret_back_tb/ret_back_synth_inst/bmg_port/ADDRA
      waveform add -signals /ret_back_tb/ret_back_synth_inst/bmg_port/DOUTA
console submit -using simulator -wait no "run"
